module VGA_Controller (
	input wire clock, clear,
	
	output wire hSync, vSync, bright
	output wire [9:0] hCOunt, vCount
);
	// This module controls the counters


endmodule