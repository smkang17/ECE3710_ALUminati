module topVGA();


endmodule