module VGA_Driver (
 input wire clock, clear,
 input wire [3:0] buttons,
 
 output wire [9:0] xLocation, yLocation,
 output wire slowPulse
);
	// Driver example but this is one of many we could use

endmodule